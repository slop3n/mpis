library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity fsm is
    port ( input : in  std_logic;
           clock : in  std_logic;
           reset : in  std_logic;
           output : out  std_logic);
end fsm;
 
architecture v1 of fsm is
begin
    -- TODO
end;